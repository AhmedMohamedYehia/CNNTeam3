//`timescale 1 ns / 1 ns
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 30.05.2020 14:45:51
// Design Name: 
// Module Name: SingleFilter_Conv_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module SingleFilter_Conv_tb();
reg clk;
//reg [3199:0] image;
//reg [799:0] filter;
//wire [1151:0] ConvImage;
reg [31:0] image [9:0][9:0];
reg [799:0] filter;
wire [31:0] ConvImage [5:0][5:0];
initial begin 
clk =0;
//these numbers are 32 bit IEEE standard form 
//imageArray = 5555522222222222222222222
//filterArray = 9999933333333333333333333
//expected result = 345
image = '{'{8'h40800000,8'h40800000,8'h40800000,8'h40800000,8'h40800000},
          '{8'h40800000,8'h40800000,8'h40800000,8'h40800000,8'h40800000},
          '{8'h40800000,8'h40800000,8'h40800000,8'h40800000,8'h40800000},
          '{8'h40800000,8'h40800000,8'h40800000,8'h40800000,8'h40800000},
          '{8'h40800000,8'h40800000,8'h40800000,8'h40800000,8'h40800000}
            };
//image=3200'h40800000408000004080000040800000408000004080000040800000408000004080000040800000408000004080000040800000408000004080000040800000408000004080000040800000408000004080000040800000404000004040000040400000404000004040000040400000408000004080000040800000408000004040000040400000404000004040000040400000404000004080000040800000408000004080000040400000404000004040000040400000404000004040000040800000408000004080000040800000404000004040000040400000404000004040000040400000408000004080000040800000408000004040000040400000404000004040000040400000404000004080000040800000408000004080000040400000404000004040000040400000404000004040000040800000408000004080000040800000408000004080000040800000408000004080000040800000408000004080000040800000408000004080000040800000408000004080000040800000408000004080000040800000;
filter=800'h3F8000003F8000003F8000003F8000003F8000003F8000003F8000003F8000003F8000003F8000003F8000003F8000003F8000003F8000003F8000003F8000003F8000003F8000003F8000003F8000003F8000003F8000003F8000003F8000003F800000;
end

always
begin 

#5 clk =~clk;
end


SingleFilter_Conv SingleLayer(clk,image,filter,ConvImage);

endmodule
